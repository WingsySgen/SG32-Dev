`define UART_MASTER_SYSCLK 1.25e+07
`define UART_BAUD_RATE 115200
`define EBR_BASED
